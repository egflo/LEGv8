`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10/20/2020 03:50:02 PM
// Design Name: 
// Module Name: instruction_memory
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module instruction_memory(PCOut, InstructionOut);

input [63:0] PCOut;
output [31:0] InstructionOut;
reg [7:0] IM[0:255];

//PC + 4 Bytes -> 1 Byte = 8 Bits -> 8 x 4 = 32 Bits

initial 
begin


/**
STORE 

------------------------------------------------------
| Opcode | Displacement | 00 | Rn(Base) | Rt (Dest)  |
------------------------------------------ ----------|
|   11   |     9        | 2  |     5    |     5      |
-----------------------------------------------------
Load/store instructions
 Rn: base register
 Displacement: constant offset from contents of base register (+/- 32
doublewords)
 Rt: destination (load) or source (store) register number
**/

/**
CBZ

-----------------------------------------
| Opcode | Relative Offset | Rt (SRC)  |
-----------------------------------------
|   8    |     19           | 5         |
----------------------------------------
**/


/**
0000 AND A & B -> ALU_Op: 1x Opcode_feild: 10001010000
0001 OR A  B -> 1x 10101010000
0010 ADD A + B -> 1x 10001011000
0110 SUBTRACT A - B ->  1x 11001011000
0111 PASS INPUT B B -> x1 xxxxxxxxxxx
1100 NOR ~ (A|B) -> 00 xxxxxxxxxxx

------------------------------------------------------
| Opcode | Src reg 2 | Shamt | Src reg 1 | Dest reg  |
------------------------------------------ ----------|
|   11   |     5     |   6   |     5     |     5     |
-----------------------------------------------------
**/

//OR X12,X9,X2
//10101010000000100000000100101100
IM[67] = 8'b0010_1100;
IM[66] = 8'b0000_0001;
IM[65] = 8'b0000_0010;
IM[64] = 8'b1010_1010;
//AND X8,X6,X2
//10001010000000100000000011001000
IM[63] = 8'b1100_1000;
IM[62] = 8'b0000_0000;
IM[61] = 8'b0000_0010;
IM[60] = 8'b1000_1010;
//SUB X5,X4,X2
//11001011000000100000000010000101
IM[59] = 8'b1000_0101;
IM[58] = 8'b0000_0000;
IM[57] = 8'b0000_0010;
IM[56] = 8'b1100_1011;
//ADD X2,X31,X1
//10001011000000010000001111100010
IM[55] = 8'b1110_0010;
IM[54] = 8'b0000_0011;
IM[53] = 8'b0000_0001;
IM[52] = 8'b1000_1011;

/**
LOAD 

------------------------------------------------------
| Opcode | Displacement | 00 | Rn(Base) | Rt (Dest)  |
------------------------------------------ ----------|
|   11   |     9        | 2  |     5    |     5     |
-----------------------------------------------------
**/

//11111000010_001100000_00_11111_01100 - LDUR X12, [X31, #96] 
//1111_1000 0100_0110 0000_0011 1110_1100
IM[51] = 8'b1110_1100;   
IM[50] = 8'b0000_0011;  
IM[49] = 8'b0100_0110; 
IM[48] = 8'b1111_1000; 

//11111000010_001011000_00_11111_01011 - LDUR X11, [X31, #88] 
//1111_1000 0100_0101 1000_0011 1110_1011
IM[47] = 8'b1110_1011;   
IM[46] = 8'b1000_0011;  
IM[45] = 8'b0100_0101; 
IM[44] = 8'b1111_1000; 

//11111000010_001010000_00_11111_01010 - LDUR X10, [X31, #80] 
//1111_1000 0100_0101 0000_0011 1110_1010
IM[43] = 8'b1110_1010;   
IM[42] = 8'b0000_0011;  
IM[41] = 8'b0100_0101; 
IM[40] = 8'b1111_1000; 

//11111000010_001001000_00_11111_01001 - LDUR X9, [X31, #72] 
//1111_1000 0100_0100 1000_0011 1110_1001
IM[39] = 8'b1110_1001;   
IM[38] = 8'b1000_0011;  
IM[37] = 8'b0100_0100; 
IM[36] = 8'b1111_1000; 

//11111000010_001000000_00_11111_01000 - LDUR X8, [X31, #64] 
//1111_1000 0100_0100 0000_0011 1110_1000
IM[35] = 8'b1110_1000;   
IM[34] = 8'b0000_0011;  
IM[33] = 8'b0100_0100; 
IM[32] = 8'b1111_1000; 

//11111000010_000111000_00_11111_00111 - LDUR X7, [X31, #56] 
//1111_1000 0100_0011 1000_0011 1110_0111
IM[31] = 8'b1110_0111;   
IM[30] = 8'b1000_0011;  
IM[29] = 8'b0100_0011; 
IM[28] = 8'b1111_1000; 

//11111000010_000110000_00_11111_00110 - LDUR X6, [X31, #48] 
//1111_1000 0100_0011 0000_0011 1110_0110
IM[27] = 8'b1110_0110;   
IM[26] = 8'b0000_0011;  
IM[25] = 8'b0100_0011; 
IM[24] = 8'b1111_1000; 

//11111000010_000101000_00_11111_00101 - LDUR X5, [X31, #40] 
//1111_1000 0100_0010 1000_0011 1110_0101 
IM[23] = 8'b1110_0101;   
IM[22] = 8'b1000_0011;  
IM[21] = 8'b0100_0010; 
IM[20] = 8'b1111_1000; 

//11111000010_000100000_00_11111_00100 - LDUR X4, [X31, #32] 
//1111_1000 0100_0010 0000_0011 1110_0100
IM[19] = 8'b1110_0100;   
IM[18] = 8'b0000_0011;  
IM[17] = 8'b0100_0010; 
IM[16] = 8'b1111_1000; 

//11111000010_000011000_00_11111_00011 - LDUR X3, [X31, #24] 
//1111_1000 0100_0001 1000_0011 1110_0011
IM[15] = 8'b1110_0011;   
IM[14] = 8'b1000_0011;  
IM[13] = 8'b0100_0001; 
IM[12] = 8'b1111_1000; 

//11111000010_000010000_00_11111_00010 - LDUR X2, [X31, #16] 
//1111_1000 0100_0001 0000_0011 1110_0010 
IM[11] = 8'b1110_0010;   
IM[10] = 8'b0000_0011;  
IM[9] = 8'b0100_0001; 
IM[8] = 8'b1111_1000; 

//11111000010_000001000_00_11111_00001 - LDUR X1, [X31, #8] 
//1111_1000_0100_0000_1000_0011_1110_0001
IM[7] = 8'b1110_0001;   //remember "little endian" convention, least significant byte is stored in the lower 
IM[6] = 8'b1000_0011;  //address, and the most significant byte is stored in the higher address 
IM[5] = 8'b0100_0000; 
IM[4] = 8'b1111_1000; 

//11111000010_000000000_00_11111_0000 - LDUR X0, [X31, #0]  
//1111_1000 0100_0000 0000_0011 1110_0001
IM[3] = 8'b1110_0000;   //remember "little endian" convention, least significant byte is stored in the lower 
IM[2] = 8'b0000_0011;  //address, and the most significant byte is stored in the higher address 
IM[1] = 8'b0100_0000; 
IM[0] = 8'b1111_1000;

end

assign InstructionOut = {IM[PCOut], IM[PCOut + 1], IM[PCOut + 2], IM[PCOut + 3]};

endmodule
